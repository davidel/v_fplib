let MAX(A, B) = ((A > B) ? A : B);
let MIN(A, B) = ((A > B) ? B : A);
let ABS(A) = (($signed(A) >= 0) ? A : -$signed(A));
let FABS(A) = ((A >= 0.0) ? A : -A);

let EXP_OFFSET(NX) = (2**(NX - 1) - 1);

// This in theory should be a typedef within the FPU interface, but then
// many HDL tools do not support hierarchical type dereferencing.
`define IEEE754(NX, NM) \
struct packed { \
  logic  sign; \
  logic [NX - 1: 0] exp; \
  logic [NM - 1: 0] mant; \
  }

